// list all paths to your design files
`include "../00_TESTBED/define.v"
`include "../01_RTL/IOTDF.v"
`include "../01_RTL/CRC.v"
`include "../01_RTL/Gray_Bin.v"
`include "../01_RTL/F_function.v"
`include "../01_RTL/Sbox.v"